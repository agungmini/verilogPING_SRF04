//untuk tampil dari binary to decimal

module bcdto7seg(in,out);

parameter bitIn= 4;
parameter bitOut= 7;

input [bitIn-1:0] in;
output [bitOut-1:0] out;

reg [bitOut-1:0] out;

always @(*)
	case(in)
		4'h0: out<= 7'b1000000;
		4'h1: out<= 7'b1111001;
		4'h2: out<= 7'b0100100;
		4'h3: out<= 7'b0110000;
		4'h4: out<= 7'b0011001;
		4'h5: out<= 7'b0010010;
		4'h6: out<= 7'b0000010;
		4'h7: out<= 7'b1111000;
		4'h8: out<= 7'b0000000;
		4'h9: out<= 7'b0010000;
		4'ha: out<= 7'b1000000;
		4'hb: out<= 7'b1000000;
		4'hc: out<= 7'b1000000;
		4'hd: out<= 7'b1000000;
		4'he: out<= 7'b1000000;
	endcase
	
endmodule
